library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity counter is
    Port ( clk : in STD_LOGIC;
           reset : in STD_LOGIC;
           count : out STD_LOGIC_VECTOR(3 downto 0));
end counter;

architecture Behavioral of counter is
    signal counter_value : unsigned(3 downto 0) := "0000";
    signal clk_divider : integer range 0 to 50000000 := 0;  -- For 50MHz clock
begin
    process(clk, reset)
    begin
        if reset = '1' then
            counter_value <= "0000";
            clk_divider <= 0;
        elsif rising_edge(clk) then
            if clk_divider = 49999999 then  -- Creates 1-second delay (50M cycles - 1)
                clk_divider <= 0;
                if counter_value = 9 then
                    counter_value <= "0000";
                else
                    counter_value <= counter_value + 1;
                end if;
            else
                clk_divider <= clk_divider + 1;
            end if;
        end if;
    end process;
    
    count <= std_logic_vector(counter_value);
    
end Behavioral;
